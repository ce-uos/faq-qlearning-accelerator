-- This file implements the Q-Learning accelerator FAQ.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use IEEE.math_real.ALL;
use IEEE.math_real.ALL;
use work.qconfig.ALL;

entity qlearning is
  Generic (
    state_width : integer := 32;
    reward_width : integer := 32;
    action_width : integer := 32;
    action_num : integer := 4;
    state_num : integer := 16;
    repsilon : integer := 80;     -- epsilon value for e-greedy
    rseed0 : integer := 12341;    -- seed for random number generator
    rseed1 : integer := 21314     -- seed for random number generator
  );
  Port ( 
    clk : in std_logic;                                        -- clock input
    enable : in std_logic;                                     -- enable input
    
    value_out : out std_logic_vector(reward_width-1 downto 0); -- value output 
    
    next_state : in std_logic_vector(state_width-1 downto 0);  -- next state generated by the environment
    state_valid : in std_logic;                                -- whether or not the state is valid
    reward : in std_logic_vector(reward_width-1 downto 0);     -- reward returned by the environment
    reward_valid : in std_logic;                               -- whether or not the reward is valid
    action : out std_logic_vector(action_width-1 downto 0);    -- action chosen in the current state
    action_valid : out std_logic                               -- whether or not the action is valid
  
  );
end qlearning;

architecture Behavioral of qlearning is

    -- some constants from the generics
    constant epsilon : unsigned(7 downto 0) := to_unsigned(repsilon, 8);
    constant seed0 : unsigned(31 downto 0) := to_unsigned(rseed0, 32);
    constant seed1 : unsigned(31 downto 0) := to_unsigned(rseed1, 32);
    
    -- learning rate shift value
    constant alpha : integer := 1;
    
    -- decay rate  shift value
    constant gamma : integer := 1;
    
    -- action write enable used for configureation with multiple action rams
    type enable_type is array (0 to action_num-1) of std_logic;
    signal awen : enable_type := (others => '0');
    
    -- these value arrray are used for the configuration wit multiple action rams
    type value_array is array (0 to action_num-1) of std_logic_vector(reward_width-1 downto 0);
    -- read action value
    signal r_avalue : value_array := (others => (others => '0'));
    -- write action value
    signal w_avalue : value_array := (others => (others => '0'));
    
    -- current action
    signal this_action : std_logic_vector(action_width-1 downto 0);
    signal this_action_valid : std_logic := '0';
    -- current value
    signal this_value : std_logic_vector(reward_width-1 downto 0);
    
    -- action chosen in the previous state
    signal last_action : std_logic_vector(action_width-1 downto 0) := (others => '0');
    signal last_action_valid : std_logic;
    -- value of the action in the previous state
    signal last_value : std_logic_vector(reward_width-1 downto 0) := (others => '0');
    -- current state
    signal state : std_logic_vector(state_width-1 downto 0);
    -- previous state
    signal last_state : std_logic_vector(state_width-1 downto 0);
    -- reward received in previous state
    signal last_reward : std_logic_vector(reward_width-1 downto 0);
    signal last_reward_valid : std_logic := '0';
    
    -- random numbers generated by LFSRs
    signal rng0 : std_logic_vector(31 downto 0);
    signal rng1 : std_logic_vector(31 downto 0);
        
    -- action rams read enable
    signal action_rams_ren : std_logic;
    -- action rams read address
    signal action_rams_ra : std_logic_vector(state_width-1 downto 0);
    -- action rams write address
    signal action_rams_wa : std_logic_vector(state_width-1 downto 0);
  
    -- registers for first pipeline stage  
    signal s1_last_reward_valid : std_logic := '0';
    signal s1_last_action : std_logic_vector(action_width-1 downto 0) := (others => '0');
    signal s1_last_value : std_logic_vector(reward_width-1 downto 0) := (others => '0');
    signal s1_last_reward : std_logic_vector(reward_width-1 downto 0);
    signal s1_qmax_value : std_logic_vector(reward_width-1 downto 0);
    signal s1_last_qmax_value : std_logic_vector(reward_width-1 downto 0);
    signal s1_last_state : std_logic_vector(state_width-1 downto 0);
    
    signal rsubv : std_logic_vector(reward_width-1 downto 0);
    signal maxvshifted : std_logic_vector(reward_width-1 downto 0);
    
    -- registers for second pipeline stage  
    signal s2_rsubv : std_logic_vector(reward_width-1 downto 0);
    signal s2_maxvshifted : std_logic_vector(reward_width-1 downto 0);
    signal s2_last_state : std_logic_vector(state_width-1 downto 0);
    signal s2_last_reward_valid : std_logic := '0';
    signal s2_last_action : std_logic_vector(action_width-1 downto 0) := (others => '0');
    signal s2_last_value : std_logic_vector(reward_width-1 downto 0) := (others => '0');
    signal s2_qmax_value : std_logic_vector(reward_width-1 downto 0);
    signal s2_last_qmax_value : std_logic_vector(reward_width-1 downto 0);
    
    -- registers for third pipeline stage 
    signal s3_last_action : std_logic_vector(action_width-1 downto 0) := (others => '0');
    signal s3_last_value : std_logic_vector(reward_width-1 downto 0) := (others => '0');
    signal s3_last_state : std_logic_vector(state_width-1 downto 0);
    signal s3_last_qmax_value : std_logic_vector(reward_width-1 downto 0);
    signal maxvshifted_plus_rsubv : std_logic_vector(reward_width-1 downto 0);
    signal s3_maxvshifted_plus_rsubv : std_logic_vector(reward_width-1 downto 0);
    signal s3_last_reward_valid : std_logic := '0';
    
    -- action and state from last pipeline stage (either 3rd or 4th)
    signal sl_last_action : std_logic_vector(action_width-1 downto 0);
    signal sl_last_state : std_logic_vector(state_width-1 downto 0);
    
    -- debug signal for the newly computed Q-value
    signal newval_dbg : std_logic_vector(reward_width-1 downto 0);
    
    -- signals for Qmax Table
    signal qmax_update : std_logic;
    signal next_qmax_read : std_logic_vector(reward_width+action_width-1 downto 0);
    signal qmax_value : std_logic_vector(reward_width-1 downto 0);
    signal qmax_action : std_logic_vector(action_width-1 downto 0);
    signal qmax_write : std_logic_vector(reward_width+action_width-1 downto 0);
    signal new_qmax : std_logic_vector(reward_width-1 downto 0);
    signal new_qmax_action : std_logic_vector(action_width-1 downto 0);
    
    signal last_qmax_value : std_logic_vector(reward_width-1 downto 0);
    signal last_qmax_action : std_logic_vector(action_width-1 downto 0);
    
    -- signals for Q-Table
    signal qtable_write : std_logic;
    signal qtable_ra : std_logic_vector(state_width+action_width-1 downto 0);
    signal qtable_wa : std_logic_vector(state_width+action_width-1 downto 0);
    signal qvalue : std_logic_vector(reward_width-1 downto 0);
    signal new_qvalue : std_logic_vector(reward_width-1 downto 0);
    
    -- signals for action generation
    signal next_random_action : std_logic_vector(action_width-1 downto 0);
    signal random_action : std_logic_vector(action_width-1 downto 0);
    signal last_random_action : std_logic_vector(action_width-1 downto 0);
    
    COMPONENT mult_24_dsps_nopipe
      PORT (
        A : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
        B : IN STD_LOGIC_VECTOR(23 DOWNTO 0);
        P : OUT STD_LOGIC_VECTOR(47 DOWNTO 0)
      );
    END COMPONENT;
    
    signal s1_qmax_value_24 : std_logic_vector(23 downto 0);
    signal s1_qmax_value_mgamma : std_logic_vector(47 downto 0);
    signal s1_qmax_value_mgamma_16 : std_logic_vector(15 downto 0);
    signal mult_gamma : std_logic_vector(23 downto 0) := X"000080"; -- 0.5
    signal s2_maxvshifted_rsubv_24 : std_logic_vector(23 downto 0);
    signal mult_alpha : std_logic_vector(23 downto 0) := X"000080"; -- 0.5
    signal s2_maxvshifted_rsubv_malpha : std_logic_vector(47 downto 0);
    signal s2_maxvshifted_rsubv_malpha_16 : std_logic_vector(15 downto 0);
begin

    gamma_mult_gen : if qconf_mult = 1 generate
        process (s1_qmax_value, last_value) begin
            if qconf_sarsa = 0 then
                s1_qmax_value_24 <= s1_qmax_value(15 downto 0) & X"00";
            else
                s1_qmax_value_24 <= last_value(15 downto 0) & X"00";
            end if;
        end process;
        
        gamma_mult : mult_24_dsps_nopipe port map (
            A => s1_qmax_value_24,
            B => mult_gamma,
            P => s1_qmax_value_mgamma
        );
        
        s1_qmax_value_mgamma_16 <= s1_qmax_value_mgamma(31 downto 16);
    end generate;
    
    alpha_mult_gen : if qconf_mult = 1 generate

        s2_maxvshifted_rsubv_24 <= std_logic_vector(signed(s2_maxvshifted) + signed(s2_rsubv)) & X"00";
        alpha_mult : mult_24_dsps_nopipe port map (
            A => s2_maxvshifted_rsubv_24,
            B => mult_alpha,
            P => s2_maxvshifted_rsubv_malpha
        );
        
        s2_maxvshifted_rsubv_malpha_16 <= s2_maxvshifted_rsubv_malpha(31 downto 16);
    end generate;

    -- instatiation of LFSRs for random number generation
    lfsr0 : entity work.lfsr_random generic map (std_logic_vector(seed0)) port map (clk, rng0);
    lfsr1 : entity work.lfsr_random generic map (std_logic_vector(seed1)) port map (clk, rng1);
    
    -- set sl_last_state and sl_last_action based on the number of pipeline stages used in the design
    stage3_last_state_action : if qconf_4stage = 0 generate
        sl_last_state <= s2_last_state;
        sl_last_action <= s2_last_action;
    end generate;
    stage4_last_state_action : if qconf_4stage = 1 generate
        sl_last_state <= s3_last_state;
        sl_last_action <= s3_last_action;
    end generate;

    -- generate one action ram per possible action
    action_rams1 : if qconf_action_rams = 1 generate
        gen_qtables : for i in 0 to action_num-1 generate
            u0 : entity work.simple_bram 
            generic map (
                memsize => state_num,
                addr_width => state_width,
                data_width => reward_width
            )
            port map (
                clk => clk,
                wen => awen(i),
                ren => state_valid,
                waddr => sl_last_state,
                raddr => next_state,
                dout => r_avalue(i),
                din => w_avalue(i)
            );
        end generate gen_qtables;
    end generate;
    
    -- generate a single RAM for the Q-table
    action_rams0 : if qconf_action_rams = 0 generate
        qtable_ra <= next_state & next_random_action;
        qtable_wa <= sl_last_state & sl_last_action;
        
        qtable : entity work.simple_bram 
        generic map (
            memsize => state_num * action_num,
            addr_width => state_width + action_width,
            data_width => reward_width
        )
        port map (
            clk => clk,
            wen => qtable_write,
            ren => '1',
            waddr => qtable_wa,
            raddr => qtable_ra,
            dout => qvalue,
            din => new_qvalue
        );
    end generate;
    
    qmax_write <= new_qmax_action & new_qmax;
    qmax_value <= next_qmax_read(reward_width-1 downto 0);
    qmax_action <= next_qmax_read((reward_width+action_width-1) downto reward_width);
    
    -- the Qmax table
    qmaxram : entity work.simple_bram
    generic map (
        memsize => state_num,
        addr_width => state_width,
        data_width => reward_width + action_width
    )
    port map (
        clk => clk,
        wen => qmax_update,
        ren => state_valid,
        waddr => sl_last_state,
        raddr => next_state,
        dout => next_qmax_read,
        din => qmax_write
    );
    
    -- Q-Learning update with 3 pipeline stages
    qlearning_update_three : if qconf_4stage = 0 generate
         process (enable, s1_last_action, s1_last_value, s1_last_reward, s1_qmax_value, s1_last_qmax_value, s1_last_reward_valid, 
                                    s2_last_action, s2_last_value, s2_rsubv, s2_maxvshifted, s2_last_reward_valid, s2_qmax_value, s2_last_qmax_value, last_value,
                                    s1_qmax_value_mgamma_16, s2_maxvshifted_rsubv_malpha_16)
            variable newval : std_logic_vector(reward_width-1 downto 0);
        begin      
            -- set some values to 0 as default
            qmax_update <= '0';
            new_qmax <= (others => '0');
            new_qmax_action <= (others => '0');
            awen <= (others => '0');
            w_avalue <= (others => (others => '0'));
            new_qvalue <= (others => '0');
            
            -- pipeline stage 1
            rsubv <= std_logic_vector(signed(s1_last_reward) - signed(s1_last_value));
            
--            if qconf_sarsa = 0 then
--                -- Q-Learning update
--                maxvshifted <= std_logic_vector(signed(s1_qmax_value) - shift_right(signed(s1_qmax_value), gamma));
--            else
--                -- SARSA update
--                maxvshifted <= std_logic_vector(signed(last_value) - shift_right(signed(last_value), gamma));
--            end if;
            
            if qconf_mult = 0 then
                if qconf_sarsa = 0 then
                    -- Q-Learning update
                    maxvshifted <= std_logic_vector(signed(s1_qmax_value) - shift_right(signed(s1_qmax_value), gamma));
                else
                    -- SARSA update
                    maxvshifted <= std_logic_vector(signed(last_value) - shift_right(signed(last_value), gamma));
                end if;
            else 
                if qconf_sarsa = 0 then
                    maxvshifted <= std_logic_vector(signed(s1_qmax_value) - signed(s1_qmax_value_mgamma_16));
                else
                    maxvshifted <= std_logic_vector(signed(last_value) - signed(s1_qmax_value_mgamma_16));
                end if;
            end if;
            
            
            -- pipeline stage 2
            if qconf_mult = 0 then
                newval := std_logic_vector(signed(s2_last_value) + signed(shift_right(signed(s2_maxvshifted) + signed(s2_rsubv), alpha)));
            else
                newval := std_logic_vector(signed(s2_last_value) + signed(s2_maxvshifted_rsubv_malpha_16));
            end if;
            newval_dbg <= newval;
            
            -- write values back to Q-table
            if qconf_action_rams = 1 then
                w_avalue(to_integer(unsigned(s2_last_action))) <= newval;
                awen(to_integer(unsigned(s2_last_action))) <= s3_last_reward_valid;
            else
                new_qvalue <= newval;
                qtable_write <= s2_last_reward_valid;
            end if;
            
            -- write max value to Qmax table
            if unsigned(newval) > unsigned(s2_last_qmax_value) then
                qmax_update <= '1';
                new_qmax <= newval;
                new_qmax_action <= s2_last_action;
            end if;
        end process;
    end generate;
    
    -- Q-Learning update with 4 pipeline stages
    qlearning_update_four : if qconf_4stage = 1 generate
        process (enable, s1_last_action, s1_last_value, s1_last_reward, s1_qmax_value, s1_last_qmax_value, s1_last_reward_valid, 
                                    s2_last_action, s2_last_value, s2_rsubv, s2_maxvshifted, s2_last_reward_valid, s2_qmax_value, s2_last_qmax_value, last_value,
                                    s3_last_action, s3_last_value, s3_maxvshifted_plus_rsubv, s3_last_reward_valid, s3_last_qmax_value,
                                    s1_qmax_value_mgamma_16, s2_maxvshifted_rsubv_malpha_16)                 
            variable newval : std_logic_vector(reward_width-1 downto 0);
        begin      
            -- set some signals to 0 as default
            qmax_update <= '0';
            new_qmax <= (others => '0');
            new_qmax_action <= (others => '0');
            awen <= (others => '0');
            w_avalue <= (others => (others => '0'));
            new_qvalue <= (others => '0');
            
            -- pipeline stage 1
            rsubv <= std_logic_vector(signed(s1_last_reward) - signed(s1_last_value));
            
            if qconf_mult = 0 then
                if qconf_sarsa = 0 then
                    -- Q-Learning update
                    maxvshifted <= std_logic_vector(signed(s1_qmax_value) - shift_right(signed(s1_qmax_value), gamma));
                else
                    -- SARSA update
                    maxvshifted <= std_logic_vector(signed(last_value) - shift_right(signed(last_value), gamma));
                end if;
            else 
                if qconf_sarsa = 0 then
                    maxvshifted <= std_logic_vector(signed(s1_qmax_value) - signed(s1_qmax_value_mgamma_16));
                else
                    maxvshifted <= std_logic_vector(signed(last_value) - signed(s1_qmax_value_mgamma_16));
                end if;
            end if;
            
            -- pipeline stage 2
            if qconf_mult = 0 then
                maxvshifted_plus_rsubv <=  std_logic_vector(shift_right(signed(s2_maxvshifted) + signed(s2_rsubv), alpha));
            else 
                maxvshifted_plus_rsubv <= s2_maxvshifted_rsubv_malpha_16;
            end if;
            
            -- pipeline stage 3
            newval := std_logic_vector(signed(s3_last_value) + signed(s3_maxvshifted_plus_rsubv));
            newval_dbg <= newval;
            
            -- write new value back to Q-table
            if qconf_action_rams = 1 then
                w_avalue(to_integer(unsigned(s3_last_action))) <= newval;
                awen(to_integer(unsigned(s3_last_action))) <= s3_last_reward_valid;
            else
                new_qvalue <= newval;
                qtable_write <= s3_last_reward_valid;
            end if;
            
            -- write max value to Qmax table
            if unsigned(newval) > unsigned(s3_last_qmax_value) then
                qmax_update <= '1';
                new_qmax <= newval;
                new_qmax_action <= s3_last_action;
            end if;
        end process;
    end generate;
    
    -- this process generates the next action based on an e-greedy policy
    epsilon_greedy_policy : if qconf_policy_random = 0 generate
        actor : process (last_value, last_action, rng0, rng1, qvalue, qmax_value, qmax_action, random_action, r_avalue) begin
            this_value <= last_value;
            this_action <= last_action;
            
            next_random_action <= rng1(action_width-1 downto 0);
            
            if unsigned(rng0(7 downto 0)) < epsilon then
                -- if random number is smaller than epsilon, use a random action
                this_action <= random_action;
                if qconf_action_rams = 1 then
                    this_value <= r_avalue(to_integer(unsigned(random_action)));
                else
                    this_value <= qvalue;
                end if;
            else
                -- if random number is larger than epsilon, use the best action
                this_action <= qmax_action;
                this_value <= qmax_value;
            end if;
        end process;
    end generate;
    
    -- this process generates the next action for the random policy
    random_policy : if qconf_policy_random = 1 generate
        actor : process (rng1, random_action, qvalue, r_avalue) begin
            next_random_action <= rng1(action_width-1 downto 0);
            
            -- use a random action as the next action
            this_action <= random_action;
            if qconf_action_rams = 1 then
                this_value <= r_avalue(to_integer(unsigned(random_action)));
            else
                this_value <= qvalue;
            end if;
        end process;
    end generate;
    
    -- this process handles internal registers, including pipeline registers
    registers : process (clk) 
    begin
        if rising_edge(clk) then
            last_value <= this_value;
            last_action <= this_action;
            this_action_valid <= state_valid;
            last_action_valid <= this_action_valid;
            state <= next_state;
            last_state <= state;
            last_reward <= reward;
            last_reward_valid <= reward_valid;
            last_qmax_value <= qmax_value;
            last_qmax_action <= qmax_action;
            random_action <= next_random_action;
            
            -- first pipeline register
            s1_last_reward_valid <= last_reward_valid;
            s1_last_action <= last_action;
            s1_last_value <= last_value;
            s1_last_reward <= last_reward;
            s1_qmax_value <= qmax_value;
            s1_last_qmax_value <= last_qmax_value;
            s1_last_state <= last_state;
            
            -- second pipeline register
            s2_last_reward_valid <= s1_last_reward_valid;
            s2_last_action <= s1_last_action;
            s2_last_state <= s1_last_state;
            s2_rsubv <= rsubv;
            s2_maxvshifted <= maxvshifted;
            s2_last_value <= s1_last_value;
            s2_qmax_value <= s1_qmax_value;
            s2_last_qmax_value <= s1_last_qmax_value;

            -- third pipeline register
            -- this is removed by vivado if the last pipeline stage is not used
            s3_last_value <= s2_last_value;
            s3_last_state <= s2_last_state;
            s3_last_action <= s2_last_action;
            s3_maxvshifted_plus_rsubv <= maxvshifted_plus_rsubv;
            s3_last_qmax_value <= s2_last_qmax_value;
            s3_last_reward_valid <= s2_last_reward_valid;
            s3_last_qmax_value <= s2_last_qmax_value;
        end if;
    end process;
    
    action <= this_action;
    action_valid <= this_action_valid;
    value_out <= this_value;

end Behavioral;
