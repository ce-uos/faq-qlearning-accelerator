library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

package qconfig is
    type logic_vector_array is array(natural range <>) of std_logic_vector(31 downto 0);
end package;
